library ieee;
use ieee.std_logic_1164.all;

entity nlui_32 is
  port (
    y   : in  std_logic_vector(31 downto 0);
    z   : out std_logic_vector(31 downto 0)
  );
end lui_32;

architecture behavioral of lui_32 is
begin

  
end behavioral;
